library verilog;
use verilog.vl_types.all;
entity SCProc_tb is
end SCProc_tb;
