module SCProcController(inst, cond_flag, rd, rs1, rs2, imm, alu_op, pc_sel, rf_wrt_data_sel, alu_in2_sel, rf_wrt_en, mem_wrt_en);
parameter INST_BIT_WIDTH = 32;
parameter REG_INDEX_BIT_WIDTH = 4;
parameter ALU_OP_WIDTH = 5;

input [INST_BIT_WIDTH - 1 : 0] inst;
input cond_flag;
output [REG_INDEX_BIT_WIDTH - 1 : 0] rd;
output [REG_INDEX_BIT_WIDTH - 1 : 0] rs1;
output [REG_INDEX_BIT_WIDTH - 1 : 0] rs2;
output [15: 0] imm;
output [ALU_OP_WIDTH - 1 : 0] alu_op;
output [1 : 0] pc_sel;
output [1 : 0] rf_wrt_data_sel;
output [1 : 0] alu_in2_sel;
output rf_wrt_en;
output mem_wrt_en;

reg [12 : 0] control_signals;
wire [8 : 0] situation;
wire [3 : 0] op;
wire [3 : 0] fn;

assign {op, fn, rd} = inst[31 : 20];
assign situation = {op, fn, cond_flag};
assign {alu_op, pc_sel, rf_wrt_data_sel, alu_in2_sel, rf_wrt_en, mem_wrt_en} = control_signals;
assign imm = inst[15 : 0];

assign rs1 = (op == 4'b0010) ? inst[23 : 20] : inst[19 : 16];
assign rs2 = (op == 4'b0011) ? inst[23 : 20] : ((op == 4'b0010) ? inst[19 : 16] : inst[15 : 12]);

always @(situation) begin
    case (situation)
9'b	110001110	: control_signals <= 13'b	0000000000010	;
9'b	110001111	: control_signals <= 13'b	0000000000010	;
9'b	110001100	: control_signals <= 13'b	0000100000010	;
9'b	110001101	: control_signals <= 13'b	0000100000010	;
9'b	110000000	: control_signals <= 13'b	0001000000010	;
9'b	110000001	: control_signals <= 13'b	0001000000010	;
9'b	110000010	: control_signals <= 13'b	0001100000010	;
9'b	110000011	: control_signals <= 13'b	0001100000010	;
9'b	110000100	: control_signals <= 13'b	0010000000010	;
9'b	110000101	: control_signals <= 13'b	0010000000010	;
9'b	110010000	: control_signals <= 13'b	0010100000010	;
9'b	110010001	: control_signals <= 13'b	0010100000010	;
9'b	110010010	: control_signals <= 13'b	0011000000010	;
9'b	110010011	: control_signals <= 13'b	0011000000010	;
9'b	110010100	: control_signals <= 13'b	0011100000010	;
9'b	110010101	: control_signals <= 13'b	0011100000010	;
9'b	010001110	: control_signals <= 13'b	0000000000110	;
9'b	010001111	: control_signals <= 13'b	0000000000110	;
9'b	010001100	: control_signals <= 13'b	0000100000110	;
9'b	010001101	: control_signals <= 13'b	0000100000110	;
9'b	010000000	: control_signals <= 13'b	0001000000110	;
9'b	010000001	: control_signals <= 13'b	0001000000110	;
9'b	010000010	: control_signals <= 13'b	0001100000110	;
9'b	010000011	: control_signals <= 13'b	0001100000110	;
9'b	010000100	: control_signals <= 13'b	0010000000110	;
9'b	010000101	: control_signals <= 13'b	0010000000110	;
9'b	010010000	: control_signals <= 13'b	0010100000110	;
9'b	010010001	: control_signals <= 13'b	0010100000110	;
9'b	010010010	: control_signals <= 13'b	0011000000110	;
9'b	010010011	: control_signals <= 13'b	0011000000110	;
9'b	010010100	: control_signals <= 13'b	0011100000110	;
9'b	010010101	: control_signals <= 13'b	0011100000110	;
9'b	010011110	: control_signals <= 13'b	1000000000110	;
9'b	010011111	: control_signals <= 13'b	1000000000110	;
9'b	011100000	: control_signals <= 13'b	0000000010110	;
9'b	011100001	: control_signals <= 13'b	0000000010110	;
9'b	001100000	: control_signals <= 13'b	0000000000101	;
9'b	001100001	: control_signals <= 13'b	0000000000101	;
9'b	110100110	: control_signals <= 13'b	0100000000010	;
9'b	110100111	: control_signals <= 13'b	0100000000010	;
9'b	110101100	: control_signals <= 13'b	0100100000010	;
9'b	110101101	: control_signals <= 13'b	0100100000010	;
9'b	110110010	: control_signals <= 13'b	0101000000010	;
9'b	110110011	: control_signals <= 13'b	0101000000010	;
9'b	110111000	: control_signals <= 13'b	0101100000010	;
9'b	110111001	: control_signals <= 13'b	0101100000010	;
9'b	110100000	: control_signals <= 13'b	0110000000010	;
9'b	110100001	: control_signals <= 13'b	0110000000010	;
9'b	110101010	: control_signals <= 13'b	0110100000010	;
9'b	110101011	: control_signals <= 13'b	0110100000010	;
9'b	110110100	: control_signals <= 13'b	0111000000010	;
9'b	110110101	: control_signals <= 13'b	0111000000010	;
9'b	110111110	: control_signals <= 13'b	0111100000010	;
9'b	110111111	: control_signals <= 13'b	0111100000010	;
9'b	010100110	: control_signals <= 13'b	0100000000110	;
9'b	010100111	: control_signals <= 13'b	0100000000110	;
9'b	010101100	: control_signals <= 13'b	0100100000110	;
9'b	010101101	: control_signals <= 13'b	0100100000110	;
9'b	010110010	: control_signals <= 13'b	0101000000110	;
9'b	010110011	: control_signals <= 13'b	0101000000110	;
9'b	010111000	: control_signals <= 13'b	0101100000110	;
9'b	010111001	: control_signals <= 13'b	0101100000110	;
9'b	010100000	: control_signals <= 13'b	0110000000110	;
9'b	010100001	: control_signals <= 13'b	0110000000110	;
9'b	010101010	: control_signals <= 13'b	0110100000110	;
9'b	010101011	: control_signals <= 13'b	0110100000110	;
9'b	010110100	: control_signals <= 13'b	0111000000110	;
9'b	010110101	: control_signals <= 13'b	0111000000110	;
9'b	010111110	: control_signals <= 13'b	0111100000110	;
9'b	010111111	: control_signals <= 13'b	0111100000110	;
9'b	001000110	: control_signals <= 13'b	0100000000000	;
9'b	001000111	: control_signals <= 13'b	0100001000000	;
9'b	001001100	: control_signals <= 13'b	0100100000000	;
9'b	001001101	: control_signals <= 13'b	0100101000000	;
9'b	001010010	: control_signals <= 13'b	0101000000000	;
9'b	001010011	: control_signals <= 13'b	0101001000000	;
9'b	001011000	: control_signals <= 13'b	0101100000000	;
9'b	001011001	: control_signals <= 13'b	0101101000000	;
9'b	001000100	: control_signals <= 13'b	0100100000000	;
9'b	001000101	: control_signals <= 13'b	0100101000000	;
9'b	001011010	: control_signals <= 13'b	0101000000000	;
9'b	001011011	: control_signals <= 13'b	0101001000000	;
9'b	001010000	: control_signals <= 13'b	0101100000000	;
9'b	001010001	: control_signals <= 13'b	0101101000000	;
9'b	001000000	: control_signals <= 13'b	0110000000000	;
9'b	001000001	: control_signals <= 13'b	0110001000000	;
9'b	001001010	: control_signals <= 13'b	0110100000000	;
9'b	001001011	: control_signals <= 13'b	0110101000000	;
9'b	001010100	: control_signals <= 13'b	0111000000000	;
9'b	001010101	: control_signals <= 13'b	0111001000000	;
9'b	001010110	: control_signals <= 13'b	0111100000000	;
9'b	001010111	: control_signals <= 13'b	0111101000000	;
9'b	001000010	: control_signals <= 13'b	0110100000000	;
9'b	001000011	: control_signals <= 13'b	0110101000000	;
9'b	001011100	: control_signals <= 13'b	0111000000000	;
9'b	001011101	: control_signals <= 13'b	0111001000000	;
9'b	001011110	: control_signals <= 13'b	0111100000000	;
9'b	001011111	: control_signals <= 13'b	0111101000000	;
9'b	011000000	: control_signals <= 13'b	0000010101010	;
9'b	011000001	: control_signals <= 13'b	0000010101010	;
        default: control_signals <= 13'b0;
    endcase
end

endmodule
